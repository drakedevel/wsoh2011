`ifdef _BUSDEC_VH
`else
`define _BUSDEC_VH 1

`define BUS_LEDS     8'h00
`define BUS_SWITCHES 8'h01
`define BUS_VGAADDR  8'h02
`define BUS_VGADATA  8'h03

`endif
