`define UC_OFFSET_JSOP_NOP 10'd1
`define UC_OFFSET_JSOP_GOTO 10'd2
`define UC_OFFSET_JSOP_IFEQ 10'd3
`define UC_OFFSET_JSOP_IFNE 10'd4
`define UC_OFFSET_JSOP_PUSH 10'd5
`define UC_OFFSET_JSOP_DUP 10'd6
`define UC_OFFSET_JSOP_DUP2 10'd7
`define UC_OFFSET_JSOP_BITOR 10'd9
`define UC_OFFSET_JSOP_BITXOR 10'd10
`define UC_OFFSET_JSOP_BITAND 10'd11
`define UC_OFFSET_JSOP_EQ 10'd12
`define UC_OFFSET_JSOP_NE 10'd13
`define UC_OFFSET_JSOP_LT 10'd14
`define UC_OFFSET_JSOP_LE 10'd15
`define UC_OFFSET_JSOP_GT 10'd16
`define UC_OFFSET_JSOP_GE 10'd17
`define UC_OFFSET_JSOP_LSH 10'd18
`define UC_OFFSET_JSOP_RSH 10'd19
`define UC_OFFSET_JSOP_URSH 10'd20
`define UC_OFFSET_JSOP_ADD 10'd21
`define UC_OFFSET_JSOP_SUB 10'd22
`define UC_OFFSET_JSOP_NOT 10'd23
`define UC_OFFSET_JSOP_BITNOT 10'd24
`define UC_OFFSET_JSOP_NEG 10'd25
`define UC_OFFSET_JSOP_VOID 10'd26
`define UC_OFFSET_JSOP_POP 10'd27
`define UC_OFFSET_OP_NOP 10'd28
`define UC_OFFSET_OP_PUSHI 10'd29
`define UC_OFFSET_OP_PUSHV 10'd30
`define UC_OFFSET_OP_BITAND 10'd31
`define UC_OFFSET_OP_GOTO 10'd32
