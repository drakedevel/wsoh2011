module cpu(/*AUTOARG*/
   // Outputs
   vgaRed, vgaGreen, vgaBlue, st__sp_2a, leds, hatch_address, Vsync,
   Hsync,
   // Inputs
   switches, rst_b, hatch_instruction, clk
   );

   /// WORLD INTERFACE ///

   /*AUTOOUTPUT*/
   // Beginning of automatic outputs (from unused autoinst outputs)
   output		Hsync;			// From Memory of cpu_memory.v
   output		Vsync;			// From Memory of cpu_memory.v
   output [31:0]	hatch_address;		// From Fetch of cpu_fetch.v
   output [7:0]		leds;			// From Memory of cpu_memory.v
   output [10:0]	st__sp_2a;		// From Decode of cpu_decode.v
   output [2:3]		vgaBlue;		// From Memory of cpu_memory.v
   output [1:3]		vgaGreen;		// From Memory of cpu_memory.v
   output [1:3]		vgaRed;			// From Memory of cpu_memory.v
   // End of automatics
   /*AUTOINPUT*/
   // Beginning of automatic inputs (from unused autoinst inputs)
   input		clk;			// To Fetch of cpu_fetch.v, ...
   input [47:0]		hatch_instruction;	// To Fetch of cpu_fetch.v, ...
   input		rst_b;			// To Fetch of cpu_fetch.v, ...
   input [7:0]		switches;		// To Memory of cpu_memory.v
   // End of automatics

   /// INTERNAL SIGNALS ///

   wire [10:0]		st__saved_sp_3a;

   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire			alu__cond_3a;		// From Execute of cpu_execute.v
   wire [4:0]		alu__op_2a;		// From Decode of cpu_decode.v
   wire [31:0]		alu__out_3a;		// From Execute of cpu_execute.v
   wire [31:0]		branch_target_4a;	// From Memory of cpu_memory.v
   wire [1:0]		c__alu_left_2a;		// From Decode of cpu_decode.v
   wire [1:0]		c__alu_right_2a;	// From Decode of cpu_decode.v
   wire [1:0]		c__branch_2a;		// From Decode of cpu_decode.v
   wire [1:0]		c__branch_3a;		// From Execute of cpu_execute.v
   wire [7:0]		c__mem_addr_3a;		// From Execute of cpu_execute.v
   wire			c__mem_write_2a;	// From Decode of cpu_decode.v
   wire			c__mem_write_3a;	// From Execute of cpu_execute.v
   wire			c__r0_2a;		// From Decode of cpu_decode.v
   wire			c__r1_2a;		// From Decode of cpu_decode.v
   wire [2:0]		c__to_push_2a;		// From Decode of cpu_decode.v
   wire [2:0]		c__to_push_3a;		// From Execute of cpu_execute.v
   wire [2:0]		c__to_push_4a;		// From Memory of cpu_memory.v
   wire [47:0]		instruction_1a;		// From Fetch of cpu_fetch.v
   wire [47:0]		instruction_2a;		// From Decode of cpu_decode.v
   wire [47:0]		instruction_3a;		// From Execute of cpu_execute.v
   wire			kill_4a;		// From Memory of cpu_memory.v
   wire [31:0]		pc_1a;			// From Fetch of cpu_fetch.v
   wire [31:0]		pc_2a;			// From Decode of cpu_decode.v
   wire [31:0]		pc_3a;			// From Execute of cpu_execute.v
   wire [31:0]		pc_4a;			// From Memory of cpu_memory.v
   wire [34:0]		r0_3a;			// From Execute of cpu_execute.v
   wire [34:0]		r1_3a;			// From Execute of cpu_execute.v
   wire			st__push_5a;		// From Writeback of cpu_writeback.v
   wire [10:0]		st__to_pop_2a;		// From Decode of cpu_decode.v
   wire [10:0]		st__to_pop_3a;		// From Execute of cpu_execute.v
   wire [10:0]		st__to_pop_4a;		// From Memory of cpu_memory.v
   wire [10:0]		st__to_pop_5a;		// From Writeback of cpu_writeback.v
   wire [34:0]		st__to_push_4a;		// From Memory of cpu_memory.v
   wire [34:0]		st__to_push_5a;		// From Writeback of cpu_writeback.v
   wire [34:0]		st__top_0_2a;		// From Decode of cpu_decode.v
   wire [34:0]		st__top_n_2a;		// From Decode of cpu_decode.v
   wire			stall_2a;		// From Decode of cpu_decode.v
   // End of automatics

   /// PIPELINE STAGES ///

   cpu_fetch Fetch(/*AUTOINST*/
		   // Outputs
		   .instruction_1a	(instruction_1a[47:0]),
		   .pc_1a		(pc_1a[31:0]),
		   .hatch_address	(hatch_address[31:0]),
		   // Inputs
		   .branch_target_4a	(branch_target_4a[31:0]),
		   .kill_4a		(kill_4a),
		   .stall_2a		(stall_2a),
		   .clk			(clk),
		   .rst_b		(rst_b),
		   .hatch_instruction	(hatch_instruction[47:0]));

   cpu_decode Decode(/*AUTOINST*/
		     // Outputs
		     .alu__op_2a	(alu__op_2a[4:0]),
		     .c__alu_left_2a	(c__alu_left_2a[1:0]),
		     .c__alu_right_2a	(c__alu_right_2a[1:0]),
		     .c__branch_2a	(c__branch_2a[1:0]),
		     .c__mem_write_2a	(c__mem_write_2a),
		     .c__to_push_2a	(c__to_push_2a[2:0]),
		     .c__r0_2a		(c__r0_2a),
		     .c__r1_2a		(c__r1_2a),
		     .instruction_2a	(instruction_2a[47:0]),
		     .pc_2a		(pc_2a[31:0]),
		     .stall_2a		(stall_2a),
		     .st__top_0_2a	(st__top_0_2a[34:0]),
		     .st__top_n_2a	(st__top_n_2a[34:0]),
		     .st__to_pop_2a	(st__to_pop_2a[10:0]),
		     .st__sp_2a		(st__sp_2a[10:0]),
		     // Inputs
		     .instruction_1a	(instruction_1a[47:0]),
		     .kill_4a		(kill_4a),
		     .pc_1a		(pc_1a[31:0]),
		     .st__push_5a	(st__push_5a),
		     .st__to_pop_5a	(st__to_pop_5a[10:0]),
		     .st__to_push_5a	(st__to_push_5a[34:0]),
		     .st__saved_sp_3a	(st__saved_sp_3a[10:0]),
		     .c__to_push_3a	(c__to_push_3a[2:0]),
		     .c__to_push_4a	(c__to_push_4a[2:0]),
		     .st__to_pop_3a	(st__to_pop_3a[10:0]),
		     .st__to_pop_4a	(st__to_pop_4a[10:0]),
		     .clk		(clk),
		     .rst_b		(rst_b));
   
   cpu_execute Execute(/*AUTOINST*/
		       // Outputs
		       .alu__cond_3a	(alu__cond_3a),
		       .alu__out_3a	(alu__out_3a[31:0]),
		       .c__branch_3a	(c__branch_3a[1:0]),
		       .c__mem_addr_3a	(c__mem_addr_3a[7:0]),
		       .c__mem_write_3a	(c__mem_write_3a),
		       .c__to_push_3a	(c__to_push_3a[2:0]),
		       .instruction_3a	(instruction_3a[47:0]),
		       .pc_3a		(pc_3a[31:0]),
		       .r0_3a		(r0_3a[34:0]),
		       .r1_3a		(r1_3a[34:0]),
		       .st__to_pop_3a	(st__to_pop_3a[10:0]),
		       // Inputs
		       .alu__op_2a	(alu__op_2a[4:0]),
		       .c__alu_left_2a	(c__alu_left_2a[1:0]),
		       .c__alu_right_2a	(c__alu_right_2a[1:0]),
		       .c__branch_2a	(c__branch_2a[1:0]),
		       .c__mem_write_2a	(c__mem_write_2a),
		       .c__to_push_2a	(c__to_push_2a[2:0]),
		       .c__r0_2a	(c__r0_2a),
		       .c__r1_2a	(c__r1_2a),
		       .instruction_2a	(instruction_2a[47:0]),
		       .kill_4a		(kill_4a),
		       .pc_2a		(pc_2a[31:0]),
		       .pc_1a		(pc_1a[31:0]),
		       .st__top_0_2a	(st__top_0_2a[34:0]),
		       .st__top_n_2a	(st__top_n_2a[34:0]),
		       .st__to_pop_2a	(st__to_pop_2a[10:0]),
		       .clk		(clk),
		       .rst_b		(rst_b));

   cpu_memory Memory(/*AUTOINST*/
		     // Outputs
		     .branch_target_4a	(branch_target_4a[31:0]),
		     .c__to_push_4a	(c__to_push_4a[2:0]),
		     .kill_4a		(kill_4a),
		     .pc_4a		(pc_4a[31:0]),
		     .st__to_pop_4a	(st__to_pop_4a[10:0]),
		     .st__to_push_4a	(st__to_push_4a[34:0]),
		     .Hsync		(Hsync),
		     .Vsync		(Vsync),
		     .leds		(leds[7:0]),
		     .vgaBlue		(vgaBlue[2:3]),
		     .vgaGreen		(vgaGreen[1:3]),
		     .vgaRed		(vgaRed[1:3]),
		     // Inputs
		     .alu__cond_3a	(alu__cond_3a),
		     .alu__out_3a	(alu__out_3a[31:0]),
		     .c__branch_3a	(c__branch_3a[1:0]),
		     .c__mem_addr_3a	(c__mem_addr_3a[7:0]),
		     .c__mem_write_3a	(c__mem_write_3a),
		     .c__to_push_3a	(c__to_push_3a[2:0]),
		     .instruction_3a	(instruction_3a[47:0]),
		     .pc_3a		(pc_3a[31:0]),
		     .r0_3a		(r0_3a[34:0]),
		     .r1_3a		(r1_3a[34:0]),
		     .st__to_pop_3a	(st__to_pop_3a[10:0]),
		     .clk		(clk),
		     .rst_b		(rst_b),
		     .switches		(switches[7:0]));

   cpu_writeback Writeback(/*AUTOINST*/
			   // Outputs
			   .st__push_5a		(st__push_5a),
			   .st__to_pop_5a	(st__to_pop_5a[10:0]),
			   .st__to_push_5a	(st__to_push_5a[34:0]),
			   // Inputs
			   .pc_4a		(pc_4a[31:0]),
			   .c__to_push_4a	(c__to_push_4a[2:0]),
			   .st__to_pop_4a	(st__to_pop_4a[10:0]),
			   .st__to_push_4a	(st__to_push_4a[34:0]),
			   .clk			(clk),
			   .rst_b		(rst_b));
   
   // synthesis translate_off
   cpu_debug Debug(/*AUTOINST*/
		   // Inputs
		   .hatch_instruction	(hatch_instruction[47:0]),
		   .kill_4a		(kill_4a),
		   .pc_1a		(pc_1a[31:0]),
		   .pc_2a		(pc_2a[31:0]),
		   .pc_3a		(pc_3a[31:0]),
		   .pc_4a		(pc_4a[31:0]),
		   .stall_2a		(stall_2a),
		   .st__push_5a		(st__push_5a),
		   .st__to_push_5a	(st__to_push_5a[34:0]),
		   .st__top_0_2a	(st__top_0_2a[34:0]),
		   .st__top_n_2a	(st__top_n_2a[34:0]),
		   .clk			(clk),
		   .rst_b		(rst_b));
   // synthesis translate_on
endmodule
